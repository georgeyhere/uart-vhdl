module uart_tx_tb();

/* TESTBENCH PARAMETERS */

/* TESTBENCH VARS */

/* DUT INSTANTIATION */

/* SIM TASKS */

/* MAIN SIM */

endmodule